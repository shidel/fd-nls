Open Watcom EXE-till-bin�r-konverterare Version 1.5
K�llkod finns tillg�nglig under Sybase Open Watcom Public License.
EXE2BIN [flaggor] exe_fil[.exe] [bin_fil]
Flaggor:
        /Q        undertryck informationsmeddelanden
        /H        visa exe-huvud
        /R        visa omlokaliseringar
        /L=<seg>  omlokalisera exe_fil till segment <seg>
        /X        ut�kat beteende, t.ex. filer > 64KB
