0.0:LABEL Version %s\n
0.1:Skapar, �ndrar eller tar bort volymetiketten f�r en disk.\n
0.2:Syntax: LABEL [enhet:][etikett] [/?]\n
0.3:  [enhet:]  Anger vilken enhet du vill s�tta etikett p�\n
0.4:  [etikett] Anger den nya etiketten du vill s�tta p� enheten\n
0.5:  /?        Visar detta hj�lpmeddelande\n
1.0:Ta bort aktuell volymetikett (Y/N)? 
1.1:Volymetikett (11 tecken, ENTER f�r ingen)? 
1.2:Volym i enhet %c saknar etikett\n
1.3:Volym i enhet %c �r %s\n
1.4:Volymens serienummer �r %04X-%04X\n
2.0:Ogiltig parameter - /%c\n
2.1:Etiketten �r f�r l�ng. Etiketten m�ste\nvara 11 tecken eller kortare..\n
2.2:Ogiltig volymetikett\n
2.3:Flera enheter angavs..\nV�lj en enhet �t g�ngen att s�tta etikett p�.\n
2.4:Ogiltig etikett\n
2.5:Inte en giltig enhet\n
2.6:Du kan inte s�tta etikett p� en n�tverksenhet\n
2.7:Du kan inte s�tta etikett p� en enhet som har\nanv�nder ASSIGN, JOIN eller SUBST.\n
2.8:Ogiltig enhet\n
