# Hj�lptext

0.0:Fria XDEL Ut�kad filborttagning   Ver
0.1:Copyright (c) 2002 Alain Mouette - GNU GPL
0.2:XDEL [/flaggor] [@][d:][s�kv�g]filnamn[.�nd]... [/flaggor]
0.3:  @             efterf�ljande filnamn �r namnet p� en fillista
0.4:  d:            enheten som xdel ska genoms�ka
0.5:  s�kv�g        katalogen d�r s�kningen ska b�rja
0.6:  filnamn.�nd   filen som ska tas bort (jokertecken till�tna)
0.7:  /D            ta bort tomma underkataloger
0.8:  /N eller /Y   ta bort angivna filer utan varning (VAR F�RSIKTIG!)
0.9:  /O            skriv �ver innan borttagning - filinneh�ll g�r F�RLORAT
0.10:  /P            fr�ga innan borttagning av varje fil
0.11:  /R            ta bort skrivskyddade filer
0.12:  /S            ta bort filer i underkataloger
0.13:  /H eller /?   detta hj�lpmeddelande
0.14:Flera filer kan anges p� kommandoraden.

# Flera meddelanden

1.0:Ta bort fil [yn]
1.1:Inget filnamn angivet
1.2:Ogiltig flagga in
1.3:Ogiltigt namn in
1.4:Kunde inte ta bort fil
1.5:Kunde inte ta bort katalog
1.6:Fel vid l�sning av fil
1.7:Fel: Slut p� minne

# Bekr�ftelse

2.0:s�kv�g
2.1:fil
2.2:�r detta vad du vill g�ra? [yn]
