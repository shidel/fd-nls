anv�ndning: BLKDROP.EXE [flaggor]

    [flaggor]      S�kert, som om du du verkligen beh�ver en flagga

BlockDrop kr�ver mus och en 386:a eller b�ttre med VGA-grafik. Jag har inte
blivit f�rdig till att l�gga till ljud �n. En dag!

Grundid�n f�r spelet �r inte j�ttekomplicerad. Beroende p� niv�n finns det ett
antal f�rglagda och speciella block slumpm�ssigt placerade i en blockstr�m.

Det finns en f�rhandsvisning av str�mmen p� den nedre h�gra delen av sk�rmen.
Den visar upp till 20 rader kommande block. N�r ett block n�r botten av
str�mmen visas det med mer detaljer ovanf�r sl�ppzonen.

Till skillnad fr�n vissa andra spel kommer block ovanf�r sl�ppzonen att falla
rakt ner och kan inte flyttas. Till slut landar de i en h�g. Fram tills att de
landar g�r de inte att interagera med.

L�t inte h�garna av block v�xa f�r h�gt. De kommer att blockera str�mmen och du
kommer att f�rlova ett liv och blir tvungen att g�ra om niv�n.

Men oroa dig inte, n�r blocken finns i h�gen s� finns det ett antal s�tt att ta
bort dem och g�ra h�gen kortare. Generellt �r det s� att en grupp av tre eller
fler block kan klickas p� och tas bort. Fler block i gruppen inneb�r fler po�ng.

Det finns h�rda block (ser lite grann ut som ett r�tt X) som inte kan klicka p�
och tas bort, oavsett hur m�nga det finns som r�r vid varandra. Du kan endast
f� bort dem genom att detonera en standardbomb i n�rheten. N�r du g�r det tas
alla block i bombens omedelbara n�rhet bort.

Det finns ocks� speciella f�rgbombsblock som kommer att ta bort alla block med
samma f�rg i h�gen. Samt andra typer av specialblock.

N�r block tas bort fr�n h�gen kommer fallande block avsiktligen att tveka lite
f�r att l�ta h�gen kollapsa fullst�ndigt innan de landar.

�h... Om du n�r en tillr�ckligt h�g niv� och r�kar se en d�skalle med korslagda
ben, klicka inte p� den. Det �r en omedelbar d�d. Det �r den enda typ av block
du aldrig vill klicka p�.

Under spelet kan du ibland anv�nda -/+ f�r att reducera eller �ka
spelhastigheten. Det har ingen effekt p� din po�ng och �r avsett f�r erfarna
spelare som kanske blir uttr�kade av de l�ngsammare niv�erna.

I b�rjan av varje niv� kan du trycka p� tabb f�r att hoppa �ver den niv�n. Men
du varnas h�rmed, niv�erna blir bara snabbare och sv�rare.

F�r n�rvarande, n�r block tas bort fr�n h�gen, kommer de endast att kollapsa
ned�t. Men jag �verv�ger att �ven l�ta dem flytta sig inn�t f�r att �ven fylla
tomma kolumner. Men jag t�nker ocks� att spelet kan blir f�r sv�rt allt f�r
snabbt. Vissa justeringar till sv�righetsgraden kan vara l�mpliga. D� kan jag,
ist�llet f�r att det bara g�r snabbare, �ka antalet samtidigt fallande block.
Men som det �r nu m�ste jag bara v�nta och se vad anv�ndarna tycker om spelet
s� h�r l�ngt.

Jag �r s�ker p� att du kan lista ut resten.

:-)
