# Language: Swedish (CP850)
# Translation by Martin Str�mberg <ams@ludd.luth.se>.
0.0:V�ntar tills anv�ndaren trycker p� en tangent
0.1:Anv�ndning
0.2:meddelande
1.0:Tryck p� en tangent f�r att forts�tta
