# Spr�k: Svenska
# Kodsida: 850
#
# �vers�ttare: Sebastian Rasmussen
#
# Blanksteg f�re text m�ste beh�llas. S�kerst�ll att inga
# blanksteg l�ggs till p� slutet av raderna.
#
0.1:\nAnv�ndning:\n
0.2:   VMSMOUNT [/H][/V|/Q|/QQ] [/L:<enh>] [/B:<str[K]>] [/LFN [/M:<n>] [/CI|/CS]]\n
0.3:   VMSMOUNT [/V|/Q|/QQ] /U\n
0.4:        /H                  - Skriver ut detta meddelande och avslutar\n
0.5:        /V                  - Utf�rlig: Skriver ut information om systemresurser\n
0.6:        /Q                  - Tystare: Utel�mnar upphovsr�ttsmeddelande\n
0.7:        /QQ                 - Tyst: Skriver inte ut n�gra meddelande alls\n
0.8:        /L:<enhetsbokstav>  - Enhetsbokstav att tilldela\n
0.9:                              (om utel�mnad, anv�nd f�rsta tillg�ngliga)\n
0.10:        /B:<storlek[K]>     - Storlek p� l�s-/skrivbuffert\n
0.11:                              (4K standard, h�gre v�rden �kar prestanda)\n
0.12:        /LFN                - L�ngt filnamnsst�d\n
0.13:        /M:<n>              - Antal manglingstecken f�r korta namn\n
0.14:                              (2 minimum, 6 maximum, 3 standard)\n
0.15:        /CI                 - K�llfilsystem �r skiftl�gesok�nsligt\n
0.16:                              (standardflagga)\n
0.17:        /CS                 - K�llfilsystem �r skiftl�gesk�nsligt\n
0.18:                              (manglar filnamn med gemena tecken)\n
0.19:        /U                  - Avinstallera\n
1.0: FEL: Enhet %c: anv�nds redan\n
1.1: FEL: Ingen enhetsbokstav tillg�nglig (LASTDRIVE �r %c)\n
1.2: FEL: DOS-version %d.%d st�ds ej. Beh�ver 5.0 eller h�gre.\n
1.3: FEL: K�r inte ovanp� VMWARE.\n
1.4: FEL: Ogiltig enhetsbokstav %c (LASTDRIVE �r %c)\n
1.5: FEL: Kan inte h�mta listan av listor!\n
1.6: FEL: Omdirigering �r inte till�ten.\n
1.7: FEL: Redan installerad. Anv�nd /U f�r att avinstallera.\n
1.8: FEL: Inga delade mappar hittade.\n
1.9: FEL: Kan inte h�mta SDA!\n
1.10: FEL: Kan inte h�mta NLS-tabellerna.\n
1.11: FEL: Buffertstorlek m�ste vara mellan %u och %u byte\n
1.12: FEL: Kan inte avinstallera.\n
1.13: FEL: Drivrutin inte installerad.\n
1.14: FEL: Manglingstecken m�ste vara mellan %u och %u\n
1.15: VARNING: TZ ogiltig eller inte definierad, tider kommer att visas i UTC.\n
1.16: VARNING: Kan inte hitta Unicode-tabell: %s
1.17: WARNING: Kan inte l�sa in Unicode-tabell: %s
1.18: WARNING: Ogiltigt filformat: %s
1.19: WARNING: Aktiv kodsida inte hittad
1.20:. Standardv�rde cp437 anv�nds\n
2.0: Monterar delade mappar i %c:\n
2.1: Framg�ngsrikt avinstallerat och borttaget fr�n minne.\n
9.0: INFO: K�r p� VMware %s Version %lu\n
9.1: INFO: UTC-skillnad �r %ld sekunder\n
9.2: INFO: Aktiv sida �r cp%d. L�ser in Unicode-tabell %s\n
9.3: INFO: Drivrutin inl�st i minne och anv�nder %u byte.\n
