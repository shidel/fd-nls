# 
#
# FreeCOM national customization file
#
#	Language: Swedish / CP850
#	Author:   Oscar Molin <oscarmolin@telia.com>
#


#  These are error messages
#
## Issued if a single character option is unknown
:TEXT_ERROR_INVALID_SWITCH
Felaktig v�xel. - /%c
.

## Issued if a longname option is unknown
:TEXT_ERROR_INVALID_LSWITCH
Felaktig v�xel. - /%s
.

## Issued if the context, the type of argument etc. is invalid
:TEXT_ERROR_ILLFORMED_OPTION
Ogiltig parameter: '%s'
.

:TEXT_ERROR_OPT_ARG
'%s' kan inte ha n�gra parametrar
.

:TEXT_ERROR_OPT_NOARG
'%s' M�ste ha en parameter
.

:TEXT_INVALID_NUMBER
Ogiltigt nummer angivet i '%s'
.

:TEXT_ERROR_CLOSE_QUOTE
Saknar omslutande citattecken: %c
.

:TEXT_ERROR_TEMPFILE
Kunde inte skapa tempor�r fil
.

:TEXT_ERROR_TOO_MANY_PARAMETERS_STR
F�r m�nga parametrar. - '%s'
.

:TEXT_ERROR_TOO_MANY_PARAMETERS
F�r m�nga parametrar.
.

:TEXT_ERROR_INVALID_PARAMETER
Felaktig parameter. - '%s'
.

:TEXT_ERROR_PATH_NOT_FOUND
S�kv�gen finns inte.
.

:TEXT_ERROR_FILE_NOT_FOUND
Kunde inte hitta filen.
.

:TEXT_ERROR_SFILE_NOT_FOUND
Kunde inte hitta filen. - '%s'
.

:TEXT_ERROR_REQ_PARAM_MISSING
Erfordrad parameter saknas.
.

:TEXT_ERROR_INVALID_DRIVE
Felaktig enhet %c:.
.

:TEXT_ERROR_BADCOMMAND#2
Felaktigt kommando eller filnamn - "%s".
.

:TEXT_ERROR_OUT_OF_MEMORY
Det finns inte tillr�ckligt med minne.
.

:TEXT_ERROR_OUT_OF_DOS_MEMORY#1
Allokering av DOS-minne misslyckades.
.

:TEXT_ERROR_CANNOTPIPE
Kan inte �ppna tempor�r fil!
.

:TEXT_ERROR_LONG_LINE_BATCHFILE
Rad #%ld i kommandofil '%s' �r f�r l�ng.
.

:TEXT_ERROR_BFILE_VANISHED
Kommandofil '%s' hittades inte.
.

:TEXT_ERROR_BFILE_LABEL
Kommandofil '%s' inneh�ller inte etiketten '%s'.
.

:TEXT_ERROR_DIRFCT_FAILED#1
%s misslyckades f�r '%s'.
.
# The next three errors must remain in this order!
:TEXT_ERROR_SET_ENV_VAR
Kunde inte ange milj�variabeln '%s'.
Milj�omr�det fullt?
.
:TEXT_ERROR_ENV_VAR_NOT_FOUND
Milj�variabeln '%s' hittades inte.
.
:TEXT_ERROR_NO_ENVIRONMENT
Inget milj�omr�de. Minnet kanske �r slut. Ange /E v�xeln.
.

# The next three errors must remain in this order!
:TEXT_ERROR_SET_ALIAS#1
Kan inte ange alias '%s'. Alias kanske �r full?
.
:TEXT_ERROR_ALIAS_NOT_FOUND#1
Alias '%s' hittades inte.
.
:TEXT_ERROR_NO_ALIAS_SEGMENT#1
Inget alias-utrymme. Minnet kan vara slut.
.

:TEXT_ERROR_SYNTAX_STR
Syntaxfel. - '%s'
.

:TEXT_ERROR_SYNTAX
Syntaxfel.
.

:TEXT_ERROR_FILENAME_TOO_LONG
Filnamnet �r f�r l�ngt. - '%s'
.

:TEXT_ERROR_SELFCOPY
Kan inte kopiera '%s' till sig sj�lv
.

:TEXT_ERROR_COMMAND_TOO_LONG
Kommandoraden f�r l�ng efter aliasut�kning!
.

:TEXT_ERROR_LINE_TOO_LONG
Raden �r f�r l�ng.  Kan inte k�ra kommando.
.

:TEXT_ERROR_HISTORY_SIZE#1
Felaktig storlek '%s'.
.

:TEXT_HISTORY_EMPTY#1
Det inga lagrade kommandon hittades.
.


:TEXT_ERROR_BAD_MCB_CHAIN
MCB kedja korrupt, eller inte FreeDOS-kompatibelt system.
.

:TEXT_ERROR_UNDEFINED_ERROR
Ok�nt fel %d.
.

:TEXT_ERROR_REGION_WARNING
Ogiltig minnesregion %d - ignoreras.
.

:TEXT_ERROR_ON_OR_OFF
ON eller OFF m�ste anges.
.

:TEXT_ERROR_BAD_VARIABLE
Felaktig variabel angiven.
.

:TEXT_ERROR_IN_MISSING#1
FOR: IN saknas.
.

:TEXT_ERROR_MISSING_PARENTHESES#1
En eller b�da parenteserna saknas.
.

:TEXT_ERROR_DO_MISSING#1
FOR: DO saknas.
.

:TEXT_ERROR_NO_COMMAND_AFTER_DO#1
FOR: Inget kommando efter DO.
.

:TEXT_ERROR_REDIRECT_FROM_FILE
Kan inte skicka indata fr�n filen '%s'.
.

:TEXT_ERROR_REDIRECT_TO_FILE
Kan inte skicka utdata till filen '%s'.
.

:TEXT_ERROR_EMPTY_REDIRECTION#1
Tom omdirigering.
.

:TEXT_ERROR_INVALID_DATE
Felaktigt datum.
.

:TEXT_ERROR_INVALID_TIME
Felaktig tid.
.

:TEXT_ERROR_NO_GOTO_LABEL
Ingen etikett angiven f�r GOTO.
.

:TEXT_CTTY_NOTIMPLEMENTED
CTTY-kommandot finns inte i denna COMMAND.COM.
.

:TEXT_ERROR_NORW_DEVICE
Felaktig eller ingen l�s/skriv-enhet '%s'.
.

:TEXT_ERROR_CTTY_DUP
Kunde inte �ndra filbeskrivning f�r TTY '%s'.
.

:TEXT_ERROR_L_NOTIMPLEMENTED
/L v�xeln �r �nnu inte implementerad.
.

:TEXT_ERROR_U_NOTIMPLEMENTED
/U v�xeln �r �nnu inte implementerad.
.

:TEXT_ERROR_WRITING_DEST
Kunde inte skriva till m�lenhet.
.

:TEXT_ERROR_CANNOT_OPEN_SOURCE
Kunde inte �ppna m�lenhet. - '%s'
.

:TEXT_ERROR_OPEN_FILE
Kunde inte �ppna filen '%s'
.

:TEXT_ERROR_READ_FILE
Kunde inte l�sa fr�n filen '%s'
.

:TEXT_ERROR_WRITE_FILE
Kunde inte skriva till filen '%s'
.

:TEXT_ERROR_LEADING_PLUS
Parametrar f�r inte b�rja med ihops�ttningstecknet '+'.
.

:TEXT_ERROR_TRAILING_PLUS
Ihops�ttningstecknet '+' f�r inte sp�ra parametrar.
.

:TEXT_ERROR_NOTHING_TO_DO
Inget att utf�ra.
.

:TEXT_ERROR_COPY
COPY misslyckades
.

:TEXT_ERROR_IF_EXIST_NO_FILENAME#1
IF EXIST: filnamn saknas
.
:TEXT_ERROR_IF_ERRORLEVEL_NO_NUMBER#1
IF ERRORLEVEL: nummer saknas
.
:TEXT_ERROR_IF_ERRORLEVEL_INVALID_NUMBER#1
IF ERRORLEVEL: ogiltigt nummer
.
:TEXT_ERROR_IF_MISSING_COMMAND#1
IF: Kommando saknas
.

:TEXT_NOT_IMPLEMENTED_YET
F�rl�t oss...inte implementerat �n.
.

:TEXT_FAILED_LOAD_STRINGS
Kunde inte ladda meddelanden i minnet.
.

:TEXT_MSG_NOTIMPLEMENTED
V�xeln /MSG har exkluderats fr�n COMMAND.COM.
.

:TEXT_MSG_ITEMS_DISPLAYED#1
%u objekt visas.
.

:TEXT_CORRUPT_COMMAND_LINE
Korrupt kommandorad. 
Detta �r ett internt fel som �r relaterat till det system som COMMAND.COM k�rs i. 
Var god rapportera detta fel.
.

:TEXT_QUOTED_C_OR_K#1
V�xlarna /C och /K f�r inte omslutas av citattecken, de ignorerades.
.

:TEXT_INIT_FULLY_QUALIFIED#1
S�kv�gen f�r COMMAND.COM m�ste vara fullst�ndig!
Det betyder att den ska inneh�lla enhetsbokstav och b�rja med ett bak�tsnedstreck.
Till exempel: C:\\FDOS

COMMAND.COM antar nu denna s�kv�g:
%s
.

:TEXT_ERROR_RESTORE_SESSION
Sessions-informationen kunde inte �terst�llas, alla lokala inst�llningar 
har g�tt f�rlorade. Se felmeddelanden ovan f�r anledningen till detta problem.
.

:TEXT_ERROR_SAVE_SESSION
Aktuell information kan inte sparas n�r programmet anv�nds. 
Se felmeddelanden ovan f�r anledningen till detta problem.
.

:TEXT_ERROR_CWD_FAILED
Enhet %c: svarar inte eller det interna minnet �r slut.
.

:TEXT_ERROR_KSWAP_ALIAS_SIZE
Speglingen misslyckades: Alias allokerar f�r mycket minne.
.


:TEXT_ERROR_KSWAP_ALLOCMEM
Speglingen misslyckades: Kunde inte allokera bortre minnet.
.

:TEXT_ERROR_ALIAS_OUT_OF_MEM#1
Slut p� alias-utrymme.
.

:TEXT_ERROR_ALIAS_NO_SUCH#1
Alias finns inte: '%s'
.

:TEXT_ERROR_ALIAS_INSERT#1
Kunde inte s�tta in alias.
.

:TEXT_ALIAS_INVALID_NAME#1
Ogiltigt namn p� alias: '%s'.
.

:TEXT_ERROR_LOADING_CONTEXT#1
Kunde inte ladda Context modulen eller Critical Error-hanteraren.
.

:TEXT_ERROR_CONTEXT_OUT_OF_MEMORY#1
Context har slut p� minne.
Om felet kvarst�r kan ni f�rs�ka med att �ka n�gon intern buffer, 
som historikbufferten eller katalogstacken.
.

:TEXT_ERROR_CONTEXT_LENGTH#1
Storleken p� context %lu byte �verskrider max-sp�rren.
�ndrar storlek p� context %u byte.
.

:TEXT_ERROR_CONTEXT_ADD_STATUS#1
Kunde inte l�gga till statusinformation till context. Detta fel kan 
indikera korrupt minne eller felaktig uppskattning av minimistorleken p� context. Var god informera prefekten f�r FreeCOM p�: freecom@freedos.org
.

:TEXT_ERROR_CONTEXT_AFTER_SWAP#1
Context-informationen �r borta efter spegling. Context �terskapas men alla alias etc. har g�tt f�rlorade.
.

#
# Informational messages
#

:TEXT_MSG_PAUSE#1
Tryck p� valfri tangent f�r att forts�tta . . .\
.

:TEXT_MSG_HISTORY_SIZE
Historikbuffertens storlek �r %d byte.
.

:TEXT_MSG_DOSKEY
DOSKEY funktioner �r redan aktiverade i prompten.
.

:TEXT_MSG_ECHO_STATE
ECHO �r %s
.

:TEXT_MSG_VERIFY_STATE
VERIFY �r %s
.

:TEXT_MSG_FDDEBUG_STATE
DEBUG utmatning �r %s.
.
:TEXT_MSG_FDDEBUG_TARGET
DEBUG utmatning skrivs ut till '%s'.
.

:TEXT_MSG_BREAK_STATE
BREAK �r %s
.

:TEXT_MSG_CURRENT_DATE
Nuvarande datum �r %s
.

## The three DATE prompts MUST be in this order!
:TEXT_MSG_ENTER_DATE_AMERICAN#1
Skriv in nytt datum (mm%sdd%s[cc]yy): \
.
:TEXT_MSG_ENTER_DATE_EUROPE#1
Skriv in nytt datum (dd%smm%s[cc]yy): \
.
:TEXT_MSG_ENTER_DATE_JAPANESE#1
Skriv in nytt datum ([cc]yy%smm%sdd): \
.

:TEXT_MSG_CURRENT_TIME
Nuvarande tid �r %s
.

:TEXT_STRING_PM#1
 pm\
.
:TEXT_STRING_AM#1
 am\
.

:TEXT_MSG_ENTER_TIME#1
Skriv in ny tid: \
.

# src-file <operation> target-file
:TEXT_MSG_COPYING
%s %s %s
.

# This prompt MUST include the pseudo key CBREAK!
# Note: This prompt ignores DOS NLS intentionally in order to
# keep interactive prompt & user-interaction in sync.
# Used by Delete all (Y/N) --> let ENTER default to NO
# Return value: a -> Yes; else -> No
:PROMPT_DELETE_ALL#1
JjNn{CR}{LF}{CBREAK}
aabb   b   b       b
Alla filer i '%s' kommer att tas bort!
Vill ni f�rts�tta (J/N)? \
.

# This prompt MUST include the pseudo key CBREAK!
# Note: This prompt ignores DOS NLS intentionally in order to
# keep interactive prompt & user-interaction in sync.
# Return value: a -> Yes; else -> No
:PROMPT_YES_NO#1
JjNn{LF}{CR}{CBREAK}{ESC}
aabb   a   a       b    b
 [Ja=RETUR, Ja=ESC] ? \
.

# This prompt MUST include the pseudo key CBREAK!
# Note: This prompt ignores DOS NLS intentionally in order to
# keep interactive prompt & user-interaction in sync.
# Attention: This prompt is issued via BIOS; any newline MUST be prefixed
#	by \r!
# Return value: a -> Yes; b -> No; c -> All; else -> Undefined
:PROMPT_CANCEL_BATCH#1
JaNnAaQq{LF}{CR}{CBREAK}{ESC}
aabbcccc   a   a       c    b
Ctrl+Break.\r
Avbryt kommandofil '%s' (Ja/Nej/Avbryt alla) ? \
.

# This prompt MUST include the pseudo key CBREAK!
# Note: This prompt ignores DOS NLS intentionally in order to
# keep interactive prompt & user-interaction in sync.
# Return value: a -> Yes; b -> No; c -> All; d -> Quit
:PROMPT_OVERWRITE_FILE#1
JjNnAaFf{BREAK}{ENTER}{ESC}
aabbccdd      d      a    b
Skriv �ver '%s' (Ja/Nej/Alla/Forts�tt) ? \
.

# This prompt MUST include the pseudo key CBREAK!
# Note: This prompt ignores DOS NLS intentionally in order to
# keep interactive prompt & user-interaction in sync.
# Return value: a -> Yes; b -> No; c -> All; d -> Quit
:PROMPT_DELETE_FILE#1
JjNnAaFf{BREAK}{ENTER}{ESC}
aabbccdd      d      a    b
Ta bort '%s' (Ja/Nej/Alla/Forts�tt) ? \
.

:TEXT_UNKNOWN_FILENAME#1
<<ok�nd>>\
.

:TEXT_DIRSTACK_EMPTY
Katalogstacken �r tom.
.

## Strings to construct the DIR output
:TEXT_DIR_HDR_VOLUME#1
 Volymen i enhet %c \
.
:TEXT_DIR_HDR_VOLUME_STRING
�r %s
.
:TEXT_DIR_HDR_VOLUME_NONE
saknar etikett
.
:TEXT_DIR_HDR_SERIAL_NUMBER
 Volymen har serienummer %04X-%04X
.
:TEXT_DIR_FTR_FILES#1
%10s fil(er)\
.
:TEXT_DIR_FTR_BYTES
   %12s byte
.
:TEXT_DIR_FTR_TOTAL_NUMBER
Totalt antal visade filer:
.
:TEXT_DIR_FTR_DIRS#1
%10s kat\
.
:TEXT_DIR_FTR_BYTES_FREE
 %15s byte lediga
.
:TEXT_DIR_DIRECTORY
Katalog i %s
.
:TEXT_DIR_DIRECTORY_WITH_SPACE
 Katalog i %s
.
:TEXT_DIR_LINE_FILENAME_WIDE#1
%-15s\
.
:TEXT_DIR_LINE_FILENAME_BARE
%-13s
.
:TEXT_DIR_LINE_FILENAME_SINGLE#1
%-13s\
.
:TEXT_DIR_LINE_FILENAME#1
%-8s %-3s \
.
:TEXT_DIR_LINE_SIZE_DIR#1
        <KAT> \
.
:TEXT_DIR_LINE_SIZE#1
   %10s \
.

:TEXT_FILE_COMPLATION_DISPLAY#1
%-14s\
.

:TEXT_MSG_PATH
PATH=%s
.
:TEXT_MSG_PATH_NONE#1
Ingen katalog att s�ka i.
.

## The following names MUST be in this order!
:TEXT_WEEKDAY_SHORT_NAME_SUNDAY#1
S�n\
.
:TEXT_WEEKDAY_SHORT_NAME_MONDAY#1
M�n\
.
:TEXT_WEEKDAY_SHORT_NAME_TUESDAY#1
Tis\
.
:TEXT_WEEKDAY_SHORT_NAME_WEDNSDAY#1
Ons\
.
:TEXT_WEEKDAY_SHORT_NAME_THURSDAY#1
Tor\
.
:TEXT_WEEKDAY_SHORT_NAME_FRIDAY#1
Fre\
.
:TEXT_WEEKDAY_SHORT_NAME_SATURDAY#1
L�r\
.

# Displayed by DEL how many files were removed.
# These three strings must be kept in order!
:TEXT_MSG_DEL_CNT_FILES#1
ingen fil togs bort.
.
:TEXT_MSG_DEL_CNT_FILES_1#1
en fil togs bort.
.
:TEXT_MSG_DEL_CNT_FILES_2#1
%u filer togs bort.
.

:TEXT_MSG_SHOWCMD_INTERNAL_COMMANDS
Tillg�ngliga interna kommandon:
.

:TEXT_MSG_SHOWCMD_FEATURES

Tillg�ngliga funktioner:
.

## Displayed within "?" <-> showcmd() to enumerate the included features
## Note the trailing single space
:TEXT_SHOWCMD_FEATURE_ALIASES#1
[alias] \
.
:TEXT_SHOWCMD_FEATURE_ENHANCED_INPUT#1
[ut�kad inmatning] \
.
:TEXT_SHOWCMD_FEATURE_HISTORY#1
[historik] \
.
:TEXT_SHOWCMD_FEATURE_FILENAME_COMPLETION#1
[filnamns-komplettering] \
.
:TEXT_SHOWCMD_FEATURE_SWAP_EXEC#1
[spegling] \
.
:TEXT_SHOWCMD_FEATURE_CALL_LOGGING#1
[start-loggning] \
.
:TEXT_SHOWCMD_FEATURE_LAST_DIR#1
[f�reg�ende katalog] \
.
:TEXT_SHOWCMD_FEATURE_KERNEL_SWAP_SHELL#1
[k�rnspegling] \
.
:TEXT_SHOWCMD_FEATURE_XMS_SWAP#1
[XMS-spegling] \
.
:TEXT_SHOWCMD_DEFAULT_TO_SWAP#1
[spegling som standard] \
.
:TEXT_SHOWCMD_FEATURE_INSTALLABLE_COMMANDS#1
[kommandon att installera] \
.
:TEXT_SHOWCMD_FEATURE_NLS#1
[DOS NLS] \
.
:TEXT_SHOWCMD_FEATURE_DIRSTACK#1
[katalogstack (PUSHD)] \
.
:TEXT_SHOWCMD_FEATURE_DEBUG#1
[FreeCOM debug] \
.

:TEXT_MSG_INIT_BYPASS_AUTOEXEC#1

Tryck F8 f�r sp�rningsl�ge, eller F5 f�r att hoppa �ver %s... \
.
:TEXT_MSG_INIT_BYPASSING_AUTOEXEC
Hoppar �ver '%s'.
.

:TEXT_MSG_VER_DOS_VERSION
DOS version %u.%u
.

:TEXT_MSG_VER_EARLY_FREEDOS
FreeDOS-k�rna (bygge 1933 eller tidigare)
.

:TEXT_MSG_VER_LATER_FREEDOS
FreeDOS-k�rna version %d.%d.%d
.


:TEXT_MSG_VER_WARRANTY
Copyright (C) 1994-2001 Tim Norman och andra.

Detta program distribueras i hop om att det ska vara anv�ndbart, 
men UTAN N�GON GARANTI; utan ens p�st�dd garanti om att det PASSAR F�R ETT VISST SYFTE. Se GNU General Public License f�r mer detaljer.

Felrapporter skickas till freedos-freecom@lists.sourceforge.net.
Uppdateringar finns tillg�ngliga p� http://freedos.sourceforge.net/freecom
.

:TEXT_MSG_VER_REDISTRIBUTION
Copyright (C) 1994-2001 Tim Norman och andra.

Detta program �r fri programvara; ni kan omdistribuera den och/eller �ndra den under reglerna definierade i GNU General Public License som det publicerats av Free Software Foundation; antingen version 2 av licensen, eller om ni �nskar, den senaste.

Felrapporter skickas till freedos-freecom@lists.sourceforge.net.
Uppdateringar finns tillg�ngliga p� http://freedos.sourceforge.net/freecom
.

:TEXT_MSG_VER_DEVELOPERS

FreeDOS kommandoprompt har utvecklats av m�nga personer, se HISTORY.TXT f�r mer detaljerad information.

Nuvarande prefekt �r Steffen Kaiser mailto:freecom@freedos.org

Felrapporter skickas till freedos-freecom@lists.sourceforge.net.
Uppdateringar finns tillg�ngliga p� http://freedos.sourceforge.net/freecom
.


# Displayed when the shell is to terminate, but has been started
# with /P option <-> shell cannot exist;
# This is a crash situation, because FreeCOM won't reach this situation
# normally otherwise
# All newlines must be prefixed by \r's !
:TEXT_MSG_REBOOT_NOW#1
\r\n\r
Kommandoprompten h�ller p� att avslutas, trots att detta\r
�r f�rbjudet (vanligtvis genom att anv�nda "/P" v�xeln).\r
Ni m�ste starta om datorn, eller om prompten k�rs i en \r
multitaskingsmilj�, st�nga av processen manuellt.\r
.

# Displayed during the initialization phase of FreeCOM, if its own
# filename could not be determined.
:TEXT_MSG_FREECOM_NOT_FOUND#1
FreeCOM:s programfil hittades inte.
Ni m�ste ange fullst�ndig s�kv�g till COMMAND.COM
som f�rsta parameter i COMMAND, till exempel:
C:\\FDOS
.


:TEXT_MEMORY_ENVIRONMENT#1
Milj�segment       : max %5u byte; ledigt %5u byte
.
:TEXT_MEMORY_CONTEXT#1
Kontext-segment    : max %5u byte; ledigt %5u byte
.	
:TEXT_MEMORY_HEAP#1
Heap               : ledigt %5lu byte
.
:TEXT_MEMORY_CTXT_ALIAS#1
\tAlias            : gr�ns %5u byte, nuvarande %5u byte, %5u objekt
.
:TEXT_MEMORY_CTXT_HISTORY#1
\tHistorik         : gr�ns %5u byte, nuvarande %5u byte, %5u objekt
.
:TEXT_MEMORY_CTXT_DIRSTACK#1
\tKatalogstack     : gr�ns %5u byte, nuvarande %5u byte, %5u objekt
.
:TEXT_MEMORY_CTXT_LASTDIR#1
\tF�reg�ende kat   : anv�nt  %5u byte, %5u objekt
.
:TEXT_MEMORY_CTXT_BATCH#1
\tKommandon�stling : anv�nt  %5u byte, %5u objekt
.
:TEXT_MEMORY_CTXT_SWAPINFO#1
\tSpelingsinfo     : anv�nt  %5u byte, %5u objekt
.


## CHCP
:TEXT_ERROR_GET_CODEPAGE#1
Kunde inte h�mta kodsida fr�n systemet.
.
:TEXT_ERROR_SET_CODEPAGE#1
Kunde inte �ndra aktuellt kodsida.
.
:TEXT_DISPLAY_CODEPAGE#1
Aktuell kodsida �r %u.
Systemets kodsida �r: %u.
.

#
# Command help text
#

:TEXT_CMDHELP_ALIAS
Visar, anger eller tar bort alias.

ALIAS [variabel[=][str�ng]]

	variabel  Anger namn p� alias.
	str�ng    Anger en serie tecken som ges till alias.


ALIAS utan parametrar visar aktuella alias.
.

:TEXT_CMDHELP_BEEP
G�r ett pip-ljud.
.

:TEXT_CMDHELP_BREAK
Anger eller tar bort ut�kad CTRL+C kontroll.

BREAK [ON | OFF]

BREAK utan parametrar visar aktuellt BREAK-inst�llning.
.

:TEXT_CMDHELP_CALL#1
Anropar ett kommandofil fr�n ett annat.

CALL [/S | /N] [/Y] [enhet:][s�kv�g]filnamn [kommandofilsparametrar]

  kommandofilsparametrar   Anger kommandoradsinformation som                                             kommandofilen beh�ver.                    
  /S tvingar, /N f�rbjuder spegling av FreeCOM.
  /Y aktiverar sp�rningsl�ge under utf�randet av kommandot.
.

:TEXT_CMDHELP_CD
Visar namnet p�, eller �ndrar, aktuell katalog.

CHDIR [enhet:][s�kv�g]
CHDIR[..]
CD [enhet:][s�kv�g]
CD[..]
CD -

  ..   Anger att ni �nskar �ndra aktuell katalog moderkatalogen.
  -    Om "f�reg�ende katalog"-funktionen �r p� byts aktuell katalog ut med          f�reg�ende katalog.

CD enhet: visar vilken katalog som �r den aktuella p� angiven enhet.
CD utan parametrar visar aktuell enhet och katalog.
Se �ven: CDD
.

:TEXT_CMDHELP_CDD
Visar namnet p�, eller �ndrar, aktuell katalog och enhet.

CDD [enhet:][s�kv�g]
CDD[..]

  ..   Anger att ni �nskar �ndra aktuell katalog moderkatalogen.
  -    Om "f�reg�ende katalog"-funktionen �r p� byts aktuell katalog ut med          f�reg�ende katalog.

Om enhet: anges �ndras aktuell arbetsenhet; detta �r den enda skillnaden 
j�mf�rt mot "CHDIR".
CDD utan parametrar visar aktuell enhet och katalog.
.

:TEXT_CMDHELP_CHCP
Visar eller anger nummer f�r aktiv kodsida.

CHCP [nnn]

  nnn   Anger ett nummer f�r en kodsida.

CHCP utan parametrar visar nummer f�r aktiv kodsida.
.

:TEXT_CMDHELP_CLS
Rensar sk�rmen.

CLS
.

:TEXT_CMDHELP_COMMAND
Startar en ny kopia av FreeCOM kommandoprompt.

COMMAND [[enhet:]s�kv�g] [enhet] [/E:nnnnn] [/L:nnnn] [/U:nnn] [/P] [/MSG]
                       [/LOW] [/Y [/[C|K] kommando]]
  [enhet:]s�kv�g  Anger s�kv�g som inneh�ller COMMAND.COM.
  enhet           Anger en h�rdvaruenhet att anv�nda f�r indata och utdata.
  /E:nnnnn        Anger startstorleken p� milj�n till nnnnn byte.
                  (nnnnn b�r vara mellan 256 och 32,768).
  /L:nnnn         Anger l�ngd p� interna buffertar (kr�ver /P).
                  (nnnn b�r vara mellan 128 och 1,024).
  /U:nnn          Anger buffertl�ngd f�r indata (kr�ver /P).
                  (nnn b�r vara mellan 128 och 255).
  /P              G�r den nya kommandoprompten permanent (kan ej avslutas).
  /MSG            Lagrar alla felmeddelanden i minnet (kr�ver /P).
  /LOW            Resident data beh�lls i det l�ga minnesomr�det.
  /Y              Stegar igenom kommandofil med /C eller /K.
  /C kommando      Utf�r angivet kommando och �terg�r till programmet.
  /K kommando      Utf�r angivet kommando och forts�tter k�ra..
.

:TEXT_CMDHELP_COPY
Kopierar en eller flera filer till en annan plats

COPY [/A | /B] k�lla [/A | /B] [+ k�lla [/A | /B] [+ ...]] [m�l
  [/A | /B]] [/V] [/Y | /-Y]

  k�lla        Anger den eller de filer som ska kopieras.
  /A           Indikerar att filen �r en ASCII-textfil.
  /B           Indikerar att filen �r en bin�r fil.
  k�lla        Anger katalog och/eller filnamn f�r de nya filerna.
  /V           Verifierar att nya filer skrivs korrekt.
  /Y           Bekr�ftelse kr�vs inte f�r att skriva �ver en befintlig fil
  /-Y          Bekr�ftelse kr�vs f�r att skriva �ver en befintlig fil

V�xeln /Y kan vara f�rinst�lld i milj�variabeln COPYCMD.
Det kan �sidos�ttas med /-Y i kommandoraden

L�gg ihop filer genom att ange en enstaka fil som m�l men flera som k�lla (anv�nd jokertecken eller formatet fil1+fil2+fil3).
.

:TEXT_CMDHELP_CTTY
�ndrar den enhet som anv�nds f�r att kontrollera systemet.

CTTY enhet

  enhet   Enheten ni vill anv�nda, t ex COM1.
.

:TEXT_CMDHELP_DATE#1
Visar eller anger datum

DATE [/D] [datum]

DATE utan parametrar visar aktuellt datum och fr�gar efter ett nytt.
Tryck RETUR f�r att beh�lla samma datum.

/D hindrar DATE fr�n att bli interaktivt.
.

:TEXT_CMDHELP_DEL#2
Tar bort en eller flera filer.

DEL [enhet:][s�kv�g]filnamn [/P] [/V]
ERASE [enhet:][s�kv�g]filnamn [/P] [/V]

  [enhet:][s�kv�g]filnamn Anger fil eller filer att ta bort. 
                          Flera filer anges med jokertecken.
  /P	Kr�ver bekr�ftelse vid borttagning av fil.
  /V	Visar alla borttagna filer.
.

:TEXT_CMDHELP_DIR#4
Visar en lista med filer och underkataloger i en katalog.

DIR [enhet:][s�kv�g][filnamn] [/P] [/W] [/A[[:]attribut]]
  [/O[[:]sortorder]] [/S] [/B] [/L] [/V]

  [enhet:][s�kv�g][filnamn]
            Anger enhet, katalog och/eller filer att visa.
            (Kan vara ut�kad eller flertalig filspecifikation)
 /P         Visar en del i taget av listan, om denna inte ryms p� sk�rmen.
 /W         Visar filer och kataloger i kolumner.
 /A         Visar endast filer med angivet attribut. (standard �r /ADHSRA)
 attribut    D  Kataloger                  R  Skrivskyddade filer
             H  Dolda filer                A  Arkivklara filer
             S  Systemfiler                -  Prefix f�r inte
 /O         Ger lista enligt sortorder.
 sortorder   N  Efter namn (alfabetisk)    S  Efter storlek (minst f�rst)
             E  Efter till�gg (alfabetisk) D  Datum och tid (�ldst f�rst)
             G  Gruppera kataloger f�rst   -  Prefix f�r omv�nd ordning
             U  Osorterade		      (Standard �r /ONG)
 /S         Visar filer i angiven katalog och filerna i dess underkataloger.
 /B         Enkelt format (Ingen inledande information och sammanfattning).
 /L         Anv�nder gemener.
 /Y eller /4 Visa 4-siffriga �rtal.

V�xlar kan f�rinst�llas med milj�variabeln DIRCMD.  
�sidos�tt dessa v�xlar med - (bindestreck), till exempel /-W.
.

:TEXT_CMDHELP_DOSKEY#1
Det externa DOSKEY-verktyget finns inbyggt i FreeCOM. Anv�nd UPP- och NEDPIL
f�r att �terkalla historiken och HISTORY f�r att visa den. Anv�nd V�NSTER-
och H�GERPIL samt END och HOME f�r att navigera inom kommandoraden och
anv�nd INSERT f�r att v�xla mellan �verskrivnings- och infogningsl�ge.
Tryck TAB f�r att komplettera aktuellt ord som filnamn; tryck tv� g�nger f�r
att visa alla matchande filer.
.

:TEXT_CMDHELP_ORIGINAL_DOSKEY#1
Redigerar kommandorader, �terkallar kommandorader, och skapar makron

DOSKEY [/v�xel ...] [makronamn=[text]]

  /BUFSIZE:storlek Anger storlek p� makro- och kommandobufferten    (standard:512)
  /ECHO:ON|OFF     Anger ECHO ON/OFF i makron                       (standard:ON)
  /FILE:fil        Anger fil med lista �ver makron
  /HISTORY         Visar alla kommandon som lagrats i minnet
  /INSERT          S�tter in nya tecken i raden n�r ni skriver
  /KEYSIZE:storlek Anger storleken p� tangentbordets type-ahead-buffert (standard:15)
  /LINE:storlek    Anger maximal storlek p� radredigerings buffert  (standard:128)
  /MACROS          Visar alla DOSKey-makron
  /OVERSTRIKE      Skriver �ver gamla tecken med nya n�r ni skriver (standard)
  /REINSTALL       Installerar en ny kopia av DOSKey
  makronamn        Namnet p� makrot som skapas
  text             Kommandon som ni vill ha i makron

UPP- och NEDPIL �terkallar kommandon
            ESC tar bort aktuellt kommando
             F7 visar lagrade kommandon
         Alt+F7 tar bort lagrade kommandon
     [tecken]F8 s�ker efter kommando som b�rjar med [tecken]
             F9 v�ljer kommando med nummer
        Alt+F10 rensar alla makrodefinitioner

Specialkoder ni kan anv�nda i DOSKey makrodefinitioner:
  $T     Kommando separator: till�ter flera kommandon i samma makro
  $1-$9  kommandofilsparametrar: likv�rdiga med %1-%9 i kommandofil
  $*     Utvidgad till allt som st�r p� kommandoraden efter makrots namn
.

:TEXT_CMDHELP_ECHO
Visar meddelanden, eller styr hurvida kommandon som k�rs ska visas visas p� sk�rmen.

  ECHO [ON | OFF]
  ECHO [meddelande]

ECHO utan parametrar visar aktuell ECHO-inst�llning.
.

:TEXT_CMDHELP_EXIT
Avslutar FreeDOS kommandoprompt.

EXIT
.

:TEXT_CMDHELP_FOR
K�r angivet kommando f�r varje fil i en grupp av filer.

FOR %variabel IN (grupp) DO kommando [kommandoparametrar]

  %variabel  Anger en utbytbar parameter.
  (grupp)    Anger en eller flera filer. Jokertecken f�r anv�ndas.
  kommando   Anger kommandot som ska utf�ras f�r varje fil.
  kommandoparametrar
             Anger parametrar och/eller v�xlar f�r det angivna kommandot.

F�r att anv�nda FOR kommandot i ett kommandofil, ange %%variabel ist�llet
f�r %variabel.
.

:TEXT_CMDHELP_GOTO
Styr kommandoprompten till en rad med given etikett i ett kommandofil.

GOTO etikett

  etikett    Anger en textstr�ng som anv�nds i kommandofil som etikett.

Ni skriver etiketten f�r sig sj�lv p� en rad, med ett kolon f�re.
.

:TEXT_CMDHELP_HISTORY#1
Historikkommando.

HISTORY [storlek]

Utan "storlek" visas det aktuella inneh�llet i historikbufferten f�r
kommandoraden.
Med "storlek" s� �ndras storleken p� historikbufferten.
.

:TEXT_CMDHELP_IF
K�r ett kommando i ett kommandoprogram om ett villkor �r sant.

IF [NOT] ERRORLEVEL tal kommando
IF [NOT] str�ng1==str�ng2 kommando
IF [NOT] EXIST filnamn kommando

  NOT               Anger att kommandoprompten ska utf�ra kommandot bara 
                    om villkoret �r falskt.                   
  ERRORLEVEL tal    Anger att villkoret �r sant om det sista programmet som 
                    k�rts returnerat en slutkod som �r lika med eller st�rre 
                    �n det angivna talet.
  kommando          Anger ett kommando som ska utf�ras om villkoret har uppn�tts.
  str�ng1==str�ng2  Anger att villkoret �r sant om de angivna textstr�ngarna 
                    �r lika.
  EXIST filnamn     Anger att villkortet �r sant om det angivna filnamnet existerar.
.

:TEXT_CMDHELP_LH
Laddar ett program till det �vre minnesomr�det.

LOADHIGH [enhet:][s�kv�g]filnamn [parametrar]
LOADHIGH [/L:region1[,minstorlek1][;region2[,minstorlek2]...] [/S]]
         [enhet:][s�kv�g]filnamn [parametrar]

/L:region1[,minstorlek1][;region2[,minstorlek2]]...
            Anger de regioner av minnet dit programmet ska laddas.  
            Region1 Anger numret f�r den f�rsta minnesregionen; minstorlek1 
            anger minimistorleken, om n�gon, f�r region1.  
            Region2 and minstorlek2 anger nummer och minimistorlek
            f�r den andra regionen osv.
            Ni kan ange hur m�nga regioner ni vill.

/S          Krymper en UMB till minimal storlek medans programmet laddas.

[enhet:][s�kv�g]filnamn
            Anger plats och namn f�r programmet.
.

:TEXT_CMDHELP_LOADFIX
Laddar ett program ovanf�r de f�rsta 64K i minnet, och k�r programmet.

LOADFIX [enhet:][s�kv�g]filnamn

Anv�nd LOADFIX f�r att ladda ett program om ni har f�tt meddelandet 
"Packad fil korrupt" n�r det laddas i det l�gre minnesomr�det.
.

:TEXT_CMDHELP_MD
Skapar en katalog.

MKDIR [enhet:]s�kv�g
MD [enhet:]s�kv�g
.

:TEXT_CMDHELP_PATH
Visar eller anger de kataloger i vilka FreeCOM s�ker efter k�rbara filer.

PATH [[enhet:]s�kv�g[;...]]
PATH ;

Skriv PATH ; om ni vill rensa alla s�kv�gsinst�llningar 
och bara s�ka i den aktuella katalogen.
PATH utan parametrar visar aktuell s�kv�g.
.

:TEXT_CMDHELP_PAUSE
Avbryter bearbetningen av ett kommandoprogram och visar meddelandet:
"Tryck p� valfri tangent f�r att forts�tta..." eller valfritt eget meddelande.

PAUSE [meddelande]
.

:TEXT_CMDHELP_PROMPT
�ndrar kommandoprompten.

PROMPT [text]

  text    Best�mmer den nya promptens utseende.

Prompten kan best� av vanliga tecken och f�ljande specialtecken:

  $Q   = (lika med-tecken)
  $$   $ (dollartecken)
  $T   Aktuell tid
  $D   Aktuellt datum
  $P   Aktuell enhet och s�kv�g
  $V   FreeDOS kommandoprompts versionsnumber
  $N   Aktuell enhet
  $G   > (st�rre �n-tecken)
  $L   < (mindre �n-tecken)
  $B   | (vertikalstreck)
  $H   Backsteg (raderar f�reg�ende tecken)
  $E   Escape-tecken (ASCII-kod 27)
  $_   Vagnretur och ny rad

PROMPT utan parametrar �terst�ller promptens standardutseende.
.

:TEXT_CMDHELP_PUSHD
L�gger nuvarande katalog till katalogstacken, med valet att
�ndra nuvarande arbetskatalog.

PUSHD [[enhet:]s�kv�g]
  D�r [enhet:]s�kv�g �r en s�kv�g till det ni vill �ndra.
.

:TEXT_CMDHELP_POPD
Tar en katalog fr�n katalogstacken, och �ndras till den.

POPD [*]
  Jockertecken ('*') parametern rensar katalogstacken.
.

:TEXT_CMDHELP_DIRS
Visar inneh�llet i en katalog.

DIRS
.

:TEXT_CMDHELP_RD
Tar bort en katalog.

RMDIR [enhet:]s�kv�g
RD [enhet:]s�kv�g
.

:TEXT_CMDHELP_REM
Markerar kommentarer i ett kommandoprogram eller CONFIG.SYS.

REM [kommentar]
.

:TEXT_CMDHELP_REN
Byter namn p� en eller flera filer/kataloger.

RENAME [enhet:][s�kv�g][katalognamn1 | filnamn1] [katalognamn2 | filnamn2]
REN [enhet:][s�kv�g][katalognamn1 | filnamn1] [katalognamn2 | filnamn2]

Ni kan inte ange enhet eller s�kv�g f�r m�lfil/katalog. 
Anv�nd kommandot MOVE f�r detta syfte.
.

:TEXT_CMDHELP_SET#1
Visar, anger eller tar bort milj�variabler.

SET [/C] [/P] [variabel=[str�ng]]

  variabel  Anger milj�variabelns namn.
  str�ng    Anger en serie tecken som tilldelas variabeln

* Om ingen str�ng anges tas angiven milj�variabel bort.

SET utan parametrar visar aktuella milj�variabler.

/C tvingar SET att beh�lla information om gemener och VERSALER i variabelnamn; som standard s� omvandlas alla gemener till versaler om milj�variabeln inte redan finns, g�r den det s� beh�ller den sitt namn.

/P Fr�gar anv�ndaren efter en str�ng som sen ges till variabeln.
.

:TEXT_CMDHELP_SHIFT#1
�ndrar numreringen av de utbytbara parametrarna i kommandoprogram.

SHIFT [DOWN]

DOWN Flyttar parameter mot b�rjan (%0); annars mot slutet.
.

:TEXT_CMDHELP_TIME#1
Visar eller st�ller in systemklockan.

TIME [/T] [tid]

Skriv TIME utan parametrar f�r att visa nuvarande tidsinst�llning och fr�ga 
efter ny inst�llning.  Tryck RETUR f�r att beh�lla samma tid.

/T hindrar TIME fr�n att bli interaktiv.
.

:TEXT_CMDHELP_TRUENAME
Visar hela s�kv�gen f�r given s�kv�g.

TRUENAME [enhet:][s�kv�g][filnamn]
.

:TEXT_CMDHELP_TYPE
Visar inneh�llet i textfiler.

TYPE [enhet:][s�kv�g]filnamn
.

:TEXT_CMDHELP_VER
Visar FreeDOS kommandoprompt version och annan information.

VER [/R] [/W] [/D] [/C]

 /R         Visar k�rnversion och annan information.
 /W         FreeDOS kommandoprompt garanti.
 /D         FreeDOS kommandoprompt omdistributionsinformation.
 /C         FreeDOS kommandoprompt medhj�lpare.
.

:TEXT_CMDHELP_VERIFY
S�ger �t FreeDOS-filsystemet att verifiera att data skrivs korrekt p� disken.

VERIFY [ON | OFF]

Skriv VERIFY utan parametrar f�r att visa nuvarande VERIFY-inst�llning.
.

:TEXT_CMDHELP_FDDEBUG
Om debug (fels�kning) �r inkompilerat i FreeDOS, s� kan detta kommando
st�nga av eller sl� p� utmatning av debug-information, 
eller visa om det �r ON eller OFF.

FDDEBUG [ON | OFF | fil]

Skriv FDDEBUG utan parameter f�r att visa nuvarande inst�llningar
f�r utmatning av debug-information.
Om en fil specificeras kommer all debug-information att skickas till den filen;
utmatningen l�ggs till sist i filen, om den redan finns. De speciella
namnen "stdout" och "stderr" kan anv�ndas f�r att vidarebefordra utmatningen 
till str�mmen standard out eller standard error.
.

:TEXT_CMDHELP_VOL
Visar diskens volymetikett och serienummer, om de finns.

VOL [enhet:]
.

:TEXT_CMDHELP_QUESTION#1
Visar en lista p� kommandon och funktioner som finns tillg�ngliga i prompten.

?
?kommando [parameter]

Den f�rsta varianten visar tillg�ngliga interna kommandon och funktioner.
Den andra kommer fr�ga om det givna kommandot ska k�ras som om
sp�rningsl�ge vore aktiverat.

.

:TEXT_CMDHELP_WHICH
S�ker och visar den exekverbara filen f�r varje givet kommando.

WHICH {kommando}
.

:TEXT_CMDHELP_MEMORY#1
Visar det interna minnet som anv�nds av FreeCOM internt

MEMORY

.

:TEXT_ERROR_COPY_PLUS_DESTINATION#1
M�let f�r COPY f�r inte inneh�lla plus ('+') tecken.
.

:TEXT_DELETE_FILE#1
Tar bort fil "%s".
.
