Detta �r hj�lpfilen f�r MORE:

MORE: Visa inneh�llet i en textfil en sk�rm �t g�ngen
  Detta program �r fri programvara, och du f�r g�rna distribuera 
  det under GNU GPL; se filen COPYING f�r vidare information.

Anv�ndning:
  kommando � MORE
  MORE fil..
  MORE < fil

Tillg�ngliga tangenter (n�r en fil visas):
  N n = N�sta fil
  Q q = Avsluta program
