	0,0: hej allesammans\n

	1,0:KITTENC - KITTEN-kompilator\n
	1,1:anv�ndning\n
	1,2:KITTENC program.exe ATTACH NLS\\program.??\n
	1,3:KITTENC program.exe ATTACH NLS\\program.DE\n
	1,4:KITTENC program.exe ATTACH NLS\\program.DE NLS\\program.fr\n
	1,5:KITTENC program.exe INFO     : visa information om spr�kresurser\n
	1,6:KITTENC program.exe DUMP     : skapa spr�kresurser\n
	1,7:KITTENC program.exe TRUNCATE : ta bort bifogade resurser\n


	2,1:filnamn <%s> kan inte �ppnas. eftersom <%s>\n
	2,2:%s: ingen s�dan fil\n
