VERSION=%0 (version %1)
LICENSE=3-klausulers BSD-licens
COPYRIGHT=Copyright (c) %1, %0
RIGHTS=Alla r�ttigheter f�rbeh�llna.

; If you want credit for your translation shown in the program, simply
; edit the LANGUAGE field and fill in the TRANSLATOR field. :-)

LANGUAGE=Svenska
TRANSLATOR=Sebastian Rasmussen

THANKS=Speciellt tack till %0 f�r �vers�ttning till %1.

LOADING=L�ser in %0...
STANDBY=V�nta, behandlar...

; The error messages in ImgView are the same as ImgEdit. There are just fewer.
; You can copy past them from ImgEdit the additional error messages will not
; hurt anything.

ERROR.VIDEO=kan inte hitta n�gon l�mplig grafikdrivrutin

ERROR.DRIVER.FIND=kan inte hitta %0-drivrutin
ERROR.DRIVER.INIT=kan inte initiera %0-drivrutin
ERROR.DRIVER.MODE=�ppnar grafikdrivrutin %0 l�ge %1

ERROR.NOHELP=hj�lp inte tillg�nlig
ERROR.FORMAT=kunde inte identifiera format f�r fil %0

ERROR.TOOBIG=bild �verskrider storleksbegr�nsning om %0 x %1 bildpunkter

ERROR.1=Ogiltig funktion
ERROR.2=Fil hittades ej
ERROR.3=S�kv�g hittades ej
ERROR.8=Slut p� minne
ERROR.201=Kontroll av dataintervall
ERROR.204=Internt pekaroperationsfel
ERROR.220=Kontroll av intern datatyp
ERROR.221=Operation st�ds ej
ERROR.222=Ogiltigt filformat
ERROR.240=Initieringsfel i grafikdrivrutin
ERROR.250=Initieringsfel i ljuddrivrutin
