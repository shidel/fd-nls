#### reserved to condition for example yes, no, quit     ####
0.0:J
0.1:N
#### Space reserved to file diskcopy.c                   ####
1.0:Ogiltig enhetsspecifikation eller icke borttagningsbart media.
1.1:Fel vid l�sning av konfigurationsfil.
1.2:Ogiltig flagga:
1.3:F�r m�nga parametrar:
1.4:File �r skrivskyddad! 
1.5:kopierad till
1.6:Filen hittade ej:
1.7:File finns redan!
1.8:Mata in K�LL-diskett i enhet
1.9:Tryck p� valfri tangent f�r att forts�tta . . .
1.10:Disk ej redo!
1.11:Kan inte �ppna avbildningsfil.
1.12:Inte tillr�ckligt med diskutrymme p� m�lenhet!
1.13:Fel vid �tkomst av avbildningsfil:
1.14:Otillr�ckligt minne f�r diskkopiering.
1.15:Anv�nder
1.16:tempor�rfil.
1.17:L�ser K�LL-diskett. . .
1.18:Mediafel vid l�sning fr�n sektor
1.19:Skriver till avbildningsfil.
1.20:Ov�ntat minnesfil.
1.21:Mata in M�L-diskett i enhet
1.22:Diskett har inte samma kapacitet som originalet.
1.23:Placera en diskett med r�tt kapacitet i enheten
1.24:eller tryck CTRL-C f�r att avbryta.
1.25:Skriver till M�L-diskett i enhet . . .
1.26:L�ser fr�n avbildningsfil.
1.27:Mediafel vid skrivning till sektor
1.28:Vill du g�ra �nnu en kopia av denna
1.29:avbildningsfil (J/N)?
1.30:disk (J/N)?
1.31:Kopiera ytterliga en disk (J/N)?
1.32:Kan inte kopiera avbildningsfil.
1.33:Problem vid l�sning fr�n avbildningsfil.
1.34:Skapar avbildningsfil . . .
1.35:Skriver avbildningsfil . . .
1.36:Problem vid skrivning till avbildningsfil.
1.37:J�mf�relsefil i sektor
1.38:Verifierar . . .
1.39:Anv�nder verifiering
1.40:Volymens serienummer �r
1.41:Sektor 0 oskrivbar! Skrivskyddad?
#### text is "Warning: options % doesn't do anything!"   ####
2.0:Varning: flagga
2.1:g�r ingenting!
#### text is "Problem copying % to %"                    ####
3.0:Problem vid kopiering av
3.1:til
#### text is "Copying % clusters, % sectors per cluster, ####
#### % bytes per sector.\n Drive size is % bytes"        ####
4.0:Kopierar
4.1:kluster
4.2:sektorer per kluster
4.3:byte per sektor.
4.4:Relevant enhetsstorlek �r
4.5:byte.
5.0:buffert om 
5.1:byte.
#### Space reserved to file parser.c                     ####
#### Text is "Syntax error on line % in                  ####
#### configuration file"                                 ####
6.0:Syntaxfel p� rad
6.1:in configuration file
6.1:i konfigurationsfil
6.2:Semantic error in configuration file
6.2:Semantisktfel i konfigurationfil
6.3:skriv inte in mer �n ett '='
#### Don't translate the following uppercase words!      ####
6.4:Ange YES eller NO
6.5:Ange NEVER eller ALWAYS
6.6:ange RECOVERY eller NORMAL
6.7:ange FAST eller FULL
6.8:ange UPDATE eller LEAVE
#### Space reserver to file recovery.c                   ####
6.10:Mediafel vid l�sning fr�n disk, skannar om...
6.11:Ol�sbar sektor vid position
#### Space reserved to file tdrvcpy.c                    ####
7.0:Placera k�lldiskett i enhet
7.1:Placera destinationsdiskett i enhet
7.2:Tryck p� valfri tangent f�r att forts�tta...
7.3:Ogiltig specifikation av k�llenhet eller icke borttagningsbart media.
7.4:Ogiltig specifikation av destinationsenhet eller icke borttagningsbart media.
7.5:Diskett har inte samma kapacitet som originalet.
7.6:Otillr�ckligt minne.
7.7:Mediafel vid l�sning fr�n sektor
7.8:Mediafel vid skrivning till sektor
7.9:Vill du kopiera tv� andra disketter (j/n)?
8.0:Placera en diskett med r�tt kapacitet i enheten
8.1:eller
8.2:eller tryck CTRL-C f�r att avbryta.
9.0:Kopierar
9.1:kluster
9.2:sektorer per kluster
9.3:byte per sektor.
9.4:Relevant enhetsstorlek �r
9.5:byte.
9.6:Kopierar . . .
9.7:Verifierar . . .
### Place reserved for the strings in the help screen ###
9.50:Copy one diskette or image file to another diskette or image file.
9.50:Kopiera en diskett eller avbildningsfil till en annan diskett/avbildningsfil.
9.51:av
9.52:k�lla
9.53:destination
9.54:k�lla:       enhet eller avbildningsfil att kopiera fr�n.
9.55:destination: enhet eller avbildningsfil att kopiera till.
9.56:varna anv�ndaren om anv�ndar�tg�rd via ljud.
9.57:verifiera l�sningar och skrivningar.
9.58:anv�nd endast minne f�r diskkopiering.
9.59:visa minnesanv�ndning (informativt).
9.60:skriv �ver destination, om den redan finns (i fallet med en avbildningsfil).
9.61:avsluta alltid automatiskt.
9.62:f�ruts�tt att disk redan finns i enhet.
9.63:g� in i �terh�mtningsl�ge f�r disk.
9.64:utf�r snabb diskkopiering (kopiera endast fyllda sektorer).
9.65:Notera:  ett minustecken efter en flagg inaktiverar flaggan.
9.66:         Du f�r ange samma enhet som k�lla och destination.
9.67:g�r inget, inkluderad f�r MS-DOS-kompatibilitet.
9.40:fr�ga inte om m�ldisk vid kopiering av avbildningsfil till samma disk.
