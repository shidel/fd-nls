FLASHROM

FLASHROM �r ett universellt verktyg f�r att s�kerhetskopiera och uppdatera
ditt system BIOS. Var f�rsiktigt vid anv�ndning d� det kan skada ditt system.
