0.0:Avg�r k�rtiden f�r ett program
0.1:Anv�ndning
1.0:K�rtiden var %f sekunder
2.0:program
