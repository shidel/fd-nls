cdrom [options]

Ett kommandoverktyg f�r inl�sning av CD/DVD-drivrutin och disktill�gg.

    [none]          F�rs�k att leta efter l�mplig drivrutin.
    search          G�r samma sak.

    help            Visa denna hj�lpsk�rm. ;)

    display         Visa f�r n�rvarande konfigurerad CD-ROM-enhet

    DRIVER_NAME     S�k inte, bara prova en specifik drivrutin.
                    (som UDVD2, GCDROM o.s.v.)

Vid s�kning, kommer den att f�rs�ka hitta och anv�nda f�ljande drivrutiner:

    AHCICD.SYS
    VIDE-CDD.SYS
    OAKCDROM.SYS
    GSCDROM.SYS
    UDVD2.SYS
    ELTORITO.SYS
    GCDROM.SYS
    UIDE.SYS

