# TEE Kitten-fil f�r SVenska
0.0:Sparar en kopia av indata till en fil och skriv ut den.
0.1:Anv�ndning
0.3:FIL(er)
0.4:L�gg till p� slutet av angiven/angivna FIL(er)
0.5:Ignorera anv�ndargenererade avbrott
0.6:Visa detta hj�lpmeddelande
1.0:Ok�nd flagga
1.1:Fel vid allokering av utrymme f�r filhandtag
1.2:Fel vid �ppning av utdatafil
1.3:Fel vid skrivning till fil
1.4:Fel vid st�ngning av fil
