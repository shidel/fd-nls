FDSHELL

FDSHELL �r en �ppenk�llkodsverion av Microsofts grafiska anv�ndargr�nssnitt DOSSHELL
Modifiera DOSSHELL.INI om det beh�vs

