# Svensk spr�kfil f�r (R)XCOPY 1.2

# fr�fr�gan och felmeddelanden
1.1:Ogiltigt antal parametrar
1.2:Ogiltigt datum
1.3:Ogiltig flagga
1.4:K�lls�kv�g f�r l�ng
1.5:Ogiltig enhetsspecifikation f�r k�lla
1.6:K�lls�kv�g hittas ej
1.7:K�lls�kv�g f�r l�ng
1.8:Destinationss�kv�g f�r l�ng
1.9:Ogiltig enhetsspecifikation f�r destination
1.10:Anger
1.11:ett filnamn
1.12:eller ett katalognamn p� m�let
1.13:Fil
1.14:Katalog
1.15:Destinationss�kv�g f�r l�ng
1.16:Kan inte utf�ra en cyklisk kopiering
1.17:Tryck p� retur f�r att forts�tta...
1.18:Fil hittades ej

# hj�lpmeddelandena
2.1:Kopierar filer och katalogtr�d.
2.2:XCOPY k�lla [destination] [/flaggor]
2.3:  k�lla        Anger katalogen och/eller namnen p� filer att kopiera.
2.4:  destination  Anger platsen och/eller namnet p� de nya filerna.
2.5:  /A           Kopierar endast filer med arkivattributet satt och �ndrar
2.6:               inte attributet.
2.7:  /C           Forts�tter kopiera �ven om fel uppst�r.
2.8:  /D[:M/D/Y]   Kopierar endast filer som har �ndrats p� eller efter det
2.9:               angivna datumet. Om inget datum anges kommer endast filer som
2.10:               �r nyare �n destinationsfilerna att kopieras.
2.11:  /E           Kopierar underkataloger, �ven om de �r tomma.
2.12:  /F           Visa fullst�ndiga k�ll- och destinationsnamn.
2.13:  /H           Kopierar g�mda och system filer s� v�l som oskyddade filer.
2.14:  /I           Om destinationen inte finns och mer �n en fil kopieras,
2.15:               f�ruts�tt att destinationen �r en katalog.
2.16:  /L           Lista filer utan att kopiera dem. (simulerar kopiering)
2.17:  /M           Kopierar endast filer med arkivattributet satt och tar bort
2.18:               akrivattributet f�r k�llfilerna efter att de kopierats.
2.19:  /N           Undertrycker fr�ga om bekr�ftelse om att du vill ta bort
2.20:               existerande destinationsfiler och hoppa �ver dessa filer.
2.21:  /P           Fr�gar om bekr�ftelse innan skapande av varje destinationsfil.
2.22:  /Q           Tyst l�ge, visa inte kopierade filnamn.
2.23:  /R           Skriv �ver skrivskydddadee filer s� v�l som oskyddade filer.
2.24:  /S           Kopierar kataloger och underkataloger, f�rutom tomma.
2.25:  /T           Skapar katalogtr�d utan att kopierar filer. Tomma kataloger
2.26:               kommer inte att kopieras. F�r att kopiera dem anv�nd flaggan /E.
2.27:  /V           Verifierar varje ny fil.
2.28:  /W           V�ntar p� en knapptryckning innan start.
2.29:  /Y           Undertrycker f�rfr�gan om att bekr�fta att du vill skriva �ver
2.30:               en existerande destinationsfil coh skriv �ver dessa filer.
2.31:  /-Y          Fr�gar om bekr�ftelse att du vill skriva �ver en existerande
2.32:               destinationsfil.
2.33:Flaggan /Y eller /N kan f�rist�llas i milj�variabeln COPYCMD.
2.34:Detta kan �sidos�ttas med /-Y p� kommandoraden.
2.35:tryck p� retur f�r mer

# fler meddelanden
1.19:fil(er) kopierad(e)
1.20:Kan inte skapa katalog
1.21:Fil kan inte kopieras p� sig sj�lv
1.22:L�s�tkomst nekad
1.23:Otillr�ckligt diskutrymme i destinationss�kv�gen
1.24:Skriv�tkomst nekad
1.25:Otillr�ckligt diskutrymme i destinationss�kv�gen
1.26:Kopierar

# f�ljande tre anv�ns i shared.inc:
25.0:Kan inte �ppna k�llfil
25.1:Kan inte skapa destination
25.2:Skrivfel vid destination

# fler bekr�ftelsemeddelanden, m�ste b�rja med versal,
# 3.2 till 3.5 m�ste alla inledas olika:
3.1:Skriv �ver
3.2:Ja
3.3:Nej
3.4:Skriv �ver alla
3.5:Hoppa �ver alla

