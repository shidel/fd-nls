# Language: Swedish (CP850)
# Translation courtesy of Martin Str�mberg <ams@ludd.luth.se>.
# Translation updated by Sebastian Rasmussen <sebras@gmail.com>.
#### Help        ####
1.0:J�mf�r tv� filer eller set av filer och visar skillnaderna mellan dem
1.1:FC [optioner] [drive1:][path1]filnamn1 [drive2][path2]filnamn2 [optioner]
1.2: /A    Visar bara den f�rsta och den sista raden f�r varje set av skillnader
1.3: /B    G�r en bin�r j�mf�relse
1.4: /C    Hantera gemener som versaler (problem med �, � och �)
1.5: /L    J�mf�r filerna som ASCII-text.
1.6: /Mn   S�tt maximal antal skillnader vid bin�r j�mf�relse till n byte.
1.7:       (default = %d, 0 = ingen begr�nsning, /M = /M0)
1.8: /N    Visa radnumren vid textj�mf�relse
1.9: /S    Ut�ka j�mf�relsen till filerna i underkatalogerna
1.10: /T    Expandera inte tabbar till mellanslag
1.11: /W    Packa tabbar och mellanslag vid textj�mf�relse
1.12: /X    Visa inte kontextrader vid textj�mf�relse
1.13: /LBn  S�tter maximalt antal konsekutiva olika ASCII-rader till n
1.14: /nnn  S�tt minsta antal konsekutiva matchande rader till nnn
1.15:       f�r omsynkronisering vid j�mf�relse
1.16: /R    Visa en kort slutrapport (alltid aktiv n�r /S anv�nds)
1.17: /Q    Visa inte listan �ver skillnader
1.18: /U    Visa filnamnen f�r filer som inte har n�gon motsvarighet
#### Messages    ####
2.0:Ogiltig option: %s
2.1:F�r m�nga filnamn
2.2:Ogiltigt filnamn
2.3:Ingen fil specificerad
2.4:Varning: filerna �r olika stora!
2.5:J�mf�relsen avslutad efter %d feltr�ffar
2.6:Inga skillnader
2.7:Varning: j�mf�relsen avbruten efter %d rader
2.8:Otillr�ckligt med minne
2.9:Fel vid �ppnande av fil %s
2.10:J�mf�r %s och %s
2.11:Ingen s�dan fil eller katalog
2.12:Omsynkronisering misslyckades: filerna �r allt f�r olika
2.13:Filerna �r olika stora
2.14:Filerna �r olika
2.15:Fil %s har ingen motsvarighet(%s)
#### Report text ####
3.0:J�mf�rde %d filer
3.1: i %d kataloger
3.2:%d filer matchar, %d filer skiljer sig
3.3:%d filer har ingen motsvarighet
