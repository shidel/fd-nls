AUTO_DONE=Behandling av uppstartsfiler klar /fCyan %1 /a7 och /fCyan %a /a7
AUTO_HELP=Skriv /fWhite %1 /fGray f�r att f� hj�lp med kommandon och navigering.
AUTO_WELCOME=V�kommentill operatigsystemet /fGreen %1 /fCyan %2 /fGray ( /s- /fYellow "%3" /fGray )
