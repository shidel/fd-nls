FDTUI

Textgr�nssnittsskal f�r FreeDOS

Copyright (C) 2017-2021 Ercan Ersoy
Detta program �r fri programvara. (GNU General Public License version 2)
                                  (GNU General Public License version 3)

Detta projekt inkluderar FDOSTUDI-biblioteket. FDOSTUI har sin egen licens.
Detta projekt inkluderar Kitten-biblioteket. Kitten har en egen licens.


Tack:

* Tack till Atnode f�r franska �vers�ttningar.
* Tack till Berki Yenig�n f�r franska �vers�ttningar.
* Tack till Eric Auer f�r Kitten-biblioteket.
* Tack till FLTK Project f�r FDOSTUI-biblioteket.
* Tack till Jerome Shidel f�r FDOSTUI-biblioteket.
* Tack till Jim Hall f�r Kitten-biblioteket.
* Tack till Mark Olesen f�r n�gra kod�ndringar och FDOSTUI-biblioteket.
* Tack till Parodper f�r spanska �vers�ttningar.
* Tack till Tom Ehlert f�r Kitten-biblioteket.
* Tack till Wilhelm Spiegl f�r tyska �vers�ttningar.


Kompilera:

  Denna programvara b�r kompileras med Open Watcom.

Bidrag:

  Om du vill bidra till detta projekt, kan du rapportera fel och g�ra
  en pull-f�rfr�ga i FDTUI-akrivet.


�ndringslogg:

* 0.7 (12-26-2021)
  * Lade till tyska �vers�ttningar.
  * Lade till spanska �vers�ttningar.
  * Uppdaterade upphovsr�ttsinformation i README.md-filen.
  * Uppdaterade tack-avsnittet i README.md-filen och README-filer.
  * Uppdaterade �ndringsloggen.

* 0.6 (12-20-2021)
  * Uppdaterade franska �ves�ttningar.
  * Uppdaterade visning av objektattribut i filhanteraren.
  * Uppdaterade hj�lpinformation.
  * Uppdaterade upphovsr�ttsinformation i README-filer.
  * Uppdaterade sk�rmbild.
  * Uppdaterade �ndringsloggen.

* 0.5 (09-20-2020)
  * Fixade n�gra typografiska fel i den franska �vers�ttningen och turkiska README.
  * Uppdaterade franska �vers�ttningar.
  * Lade till en ny franska README-fil.
  * Uppdaterade �ndringsloggen.

* 0.4 (05-28-2020)
  * �ndrade namn p� denna programvara till "FDTUI".
  * Fixade hj�lpinformation f�r lokalisering.
  * Fixade n�gra typografiska fel.
  * Uppdaterade franska �vers�ttningar.
  * Uppdaterade .gitignore-fil.
  * Tog bort attributet k�rbar f�r k�llkod.
  * Uppdaterade LICENSE, README.md, engelsk README och turkiska README-filer.
  * Tog bort fransk README-fil.
  * Uppdaterade �ndringsloggen.

* 0.3 (12-09-2018)
  * �ndrade f�rgtema.
  * �ndrade menyrad.
  * Uppdaterade spr�kfiler.
  * Tog bort on�diga rade i DOSSHELL.FR-filen.
  * Fixade "Visa arkivattribut" och fixade "Visa g�mda objekt"-kryssrutor
    i filhanteraren.
  * Inaktivera ESC-tangenten.
  * Bytade ut katalogtr�det.
  * Fixade n�gra typografiska fel.
  * Fixade fel vid val av drivrutin i listbox med tangentbord.
  * Fixade objektattribut som inte visades vid byte av enhet och fel vid
    �ppning av filhanterare.
  * Dela upp headerfiler och k�llkodsfiler.
  * Fixade hj�lpparameter.
  * �ndrade �ndelser f�r header-filer fr�n ".h" till ".hpp"
  * Ersatte sk�rmrensning som standard funktion fr�n Open Watcom ist�llet
    f�r CLS-kommando.
  * Fixade alla varningar.
  * Lade till licensinformation f�r GNU GPL version 2.
  * Uppdaterade �ndringsloggen.

* 0.2 (09-24-2018)
  * F�rgrundsf�rg f�r inaktiverade menyobjekt har �ndrats till gr�. Men den
    ser r�d ut.
  * �ndrade standardv�rden till att visa arkivobjekt och skrivskyddade objekt.
  * Lade till en paus vid avslutande kommando vid k�rning av kommando.
  * Uppdaterade engelska och turkiska �vers�ttningar.
  * Korrigerade nyradstecken anv�nda i n�gra filer ist�llet f�r felaktiga
    nyradstecken.
  * Uppdaterade �ndringsloggen.

* 0.1 (07-13-2018)
  * Skapade f�rsta versionen.


Not:

* FreeDOS �r ett varum�rke fr�n Jim Hall.
