0.0:Avg�r k�rtiden f�r ett program
1.0:K��rdtiden var %f sekunder
2.0:program
