DOSUSB

DOSUSB �r en drivrutin f�r vissa USB-styrkort med �ppen k�llkod.
F�r n�rvarande fungerar den enbart med UHCI-styrkort, d.v.s. USB 1.1
Det finns �nnu inget st�d f�r USB 2.0 och USB 3.0.
