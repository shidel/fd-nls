2.0:Ogiltig parameter\n
0.0:    SORT [/R] [/+num] [/A] [/?] [fil]\n
0.1:    /R    Omv�nd ordning\n
0.2:    /A    Anv�nd ASCII sorteringsordning ist�llet f�r den f�r COUNTRY\n
0.3:    /+num b�rja sortera med kolumn num, 1-baserat\n
0.4:    /?    hj�lp\n
2.1:Fel vid l�sning av NLS-ordningstabell\n
2.2:Anv�nd ASCII sorteringsordning (gammal DOS-version)\n
2.3:SORT: Kan inte �ppna fil '%s' f�r l�sning\n
2.5:SORT: otillr�ckligt minne\n
2.6:SORT: antal poster �verstiger maximum\n
