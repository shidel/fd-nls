Detta �r readme:n f�r FreeDOS-programmet TREE

Visar katalogstrukturen f�r en enhet eller en s�kv�g.

Anv�ndning:  TREE [/A] [/F] [S�KV�G]
  /A     Anv�nd ASCII linjeritningstecken
  /F     Visar filer i kataloger (ist�llet f�r enbart kataloger)
  S�KV�G Var katalogtr�det ska visas fr�n, standardv�rdet �r
         den aktuella katalogen.

Detta program har st�d f�r internationella tecken via biblioteket
"Cats" (catopen/catgets implementation f�r DOS).  Du kan h�mta
biblioteket "Cats" fr�n http://www.freedos.org/jhall/cats

TREE distribueras under GNU GPL.  Se filen COPYING
f�r vidare information.

