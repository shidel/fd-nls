# Language: Sveden (CP 865)
# Translated by: unknown
# Last update: unknown
2.0:Ogiltig parameter\r\n
0.0:    SORT [/R] [/+num] [/A] [/?] [fil]\r\n
0.1:    /R    Omv�nd ordning\r\n
# 0.2:    /N    Aktivera NLS-st�d\r\n - borttagen 7/2004
0.2:    /A    Anv�nd ASCII sorteringsordning ist�llet f�r den f�r COUNTRY\r\n
0.3:    /+num b�rja sortera med kolumn num, 1-baserat\r\n
0.4:    /?    hj�lp\r\n
2.1:Fel vid l�sning av NLS-ordningstabell\r\n
2.2:Anv�nd ASCII sorteringsordning (gammal DOS-version)\r\n
2.3:SORT: Kan inte �ppna fil
2.4: f�r l�sning\r\n
2.5:SORT: otillr�ckligt minne\r\n
2.6:SORT: antal poster �verstiger maximum\r\n
