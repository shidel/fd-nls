# Translation by Martin Str�mberg <ams@ludd.luth.se>
0.0:V�ntar tills anv�ndaren trycker p� en tangent fr�n en lista av val
0.1:val
0.2:text
0.3:Specificerar vilka tangenter som �r giltiga. Standardv�rde �r:
0.4:Visa inte valen efter prompten
0.5:Versaler skilda fr�n gemener
0.6:**Ignorerad, f�r kompatibilitet med MS-DOS
0.7:Texten som ska visas som prompt
0.8:Ljud en signal n�r prompten visas
3.0:jn

0.9:Felaktig tidssyntax. F�rv�ntade formen Tc,nn eller T:c,nn
0.10:Standardv�rde f�r tidsgr�ns finns ej bland angivna val (eller standardv�rde)
