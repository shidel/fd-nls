
K�llkoden f�r denna version av $OS_NAME$ och den inkluderande programvaran
�r tillg�nglig p� CD-ROM:en och USB-mediat. Den kan ocks� erh�llas via
$OS_NAME$ projektets webbplats p� $URL$
