vdelete [flaggor]

Ta bort rad p� aktuell position.

    [inga]      Ta bort rad
    n           Ta bort n rader
    /A n        S�tt textattribut till n.
    /B f�rg     S�tt textattribut f�r bakgrunden till f�rg (eller v�rde).
    /F f�rg     S�tt textattribut f�r f�rgrunden till f�rg (eller v�rde).
    /G          Global borttaning
    /L          Lokal borttaning. (Standard)
    /K n        Anv�nd n ist�llet f�r ramtecken f�r att identifiera ramar.

