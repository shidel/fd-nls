
$OS_NAME$ $OS_VERSION$ diskettutg�va 

FreeDOS-k�rnen och de flesta program i denna distribution lyder under villkoren
f�r diverse versioner av General Public License (GPL) och andra �ppenk�llkods-
licenser. F�r vidare information, bes�k FreeDOS-projektets webbplats p�
$URL$

FreeDOS �r ett varum�rke av Jim Hall, 2001-$YEAR$
