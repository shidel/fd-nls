# svedish, sv, cp 858 

99.0:Skriver ut lokaliserade meddelanden (fr�n localize.*)
99.1:Skriver ut meddelande nummer x.y eller, om inte tillg�ngligt, texten efter @@@\r\n(och slutligen ekar [et.c], om n�got)
99.2:Errorlevel: 0 om okej, 1 om ingen localize.* hittades eller inget meddelande x.y fanns inuti.
