
# Critical error national customization file
#
#	Language: Swedish / CP850
#	Author:   Oscar Molin <oscarmolin@telia.com>
# 

#
## Primary strings
S2
BLOCK_DEVICE: Fel %1 enhet %A: %2 omr�de: %3
S3
CHAR_DEVICE: Fel %1 enhet %A: %3

## kind of operation
S0
READ: l�ser fr�n
S1
WRITE: skriver till

## kind of failed area of block devices
S4
DOS: DOS
S5
FAT: FAT
S6
ROOT: Rot
S7
DATA: Data

## action strings
S8
IGNORE: (I)gnorera
S9
RETRY: (N)ytt f�rs�k
S10
ABORT: (A)vbryt
S11
FAIL: (F)orts�tt
## keys associated with the actions
S14 (compacted)
KEYS_IGNORE: iI
KEYS_RETRY:  rR
KEYS_ABORT:  aA
KEYS_FAIL:   fF
## embedded strings
S12
QUESTION:  ? %.
S13
DELIMITER: , %.

## Error strings
UNKNOWN: Ok�nd fel-kod
S15
0: f�rs�k att bryta skrivskyddet
1: ok�nd typ f�r drivrutin
2: enhet inte klar
3: drivrutin fick ok�nt kommando
4: datafel (fel CRC)
5: ogiltig strukturl�ngd p� drivrutinsbeg�ran
6: s�kfel
7: ok�nd mediatyp
8: sektorn hittades inte
9: slut p� papper i skrivaren
10: skrivfel
11: l�sfel
12: allm�nt fel
13: delningsfel
14: l�s fel
15: felaktigt diskbyte
16: FCB ej tillg�nglig
17: delningsbuffer overflow
18: codepage st�mmer inte
19: ingen input
20: otillr�ckligt diskutrymme
