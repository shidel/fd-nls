Enkel bildvisare

anv�ndning: IMGVIEW.EXE [filnamn] [filnamn] [...]

    [filnamn]       Ange fil att visa.

Endast begr�nsat st�d f�r icke-inbyggda filformat (som BMP).

Under visning...

    PgUp    F�reg�ende bild
    PgDown  N�sta bild
    Enter   Visa om
    Escape  Avsluta
