DOSUTIL

En samling anv�ndbara kommandofilsverktyg
