0.0:�vers�tter tecken
0.1:Anv�ndning:
1.0:Inte tillr�ckligt med argument
1.1:F�r m�nga argument
2.0:fil
