FLASHROM

FLASHROM is a universal tool for backing up and updating your system BIOS.
ditt system BIOS. Var f�rsiktigt vid anv�ndning d� det kan skada ditt system.
