DOSUTIL

En samling anv�ndbara BATCH-filsverktyg
