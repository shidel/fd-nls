[repository]

	Caption=FreeDOS 1.4 nedladdningar
	Description=Programvaruförråd för hämtningar och uppdateringar för FreeDOS 1.4
