0.0:Visa ett hj�lp�mne
0.1:Anv�ndning:
0.2:�mne
0.3:Milj�:
0.4:Sidvisningsprogram f�r att visa en textfil
0.5:Katalog som inneh�ller dina hj�lpfiler
0.6:F�redraget spr�k f�r dina hj�lpfiler
1.0:Kan inte k�ra sidvisningprogram.
