veach [flaggor]

G�r n�gonting f�r varje objekt i en lista.

    /S          Sl� p� list sortering.
    /L          Visa listinneh�ll.
    /F fil      L�gg till objet till lista fr�n fil.
    /I          L�gg till objekt till lista fr�n standard in.
    /D spec     L�gg till filnamn som matchar spec till listan.
    /A +/-      Modifierar /d-flaggan till att aktivera alla filer/kataloger
    /C          N�t /x-flaggan anv�ndas, till�t forts�ttning trots ett
                fel i underprocessen.
    /X [kmdrd]  K�r objekt med kommandorad och alla efterf�ljande flaggor
                skickas vidare till underprocessen. * expanderas till
		objektet, # �r antalet objekt och @ �r objektets index.
		Om ingen kommandoradsdata f�ljer p� /x-flaggan antas *.

   tba         (Fortfarande under utveckling, mer kommer att annonseras)

