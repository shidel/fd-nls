[repository]

	Caption=Senaste och instabilt
	Description=De senaste programvupaketversionerna att för att hämta eller uppdatera FreeDOS

[base]
	Caption=FreeDOS-bas
	Description=Program som tillhandahåller funktionaliteten hos klassiska DOS

[tools]
	Caption=Grundläggande verktyg
	Description=Program och verktyg som är fundamentala för FreeDOS-uppelvelsen

[apps]
	Caption=Applikationer
	Description=Interaktiva program och applikationer som är mer än bara kommandoradsverktyg

[archiver]
	Caption=Arkiverare
	Description=Verktyg för att komprimera filer och skapa arkiv

[boot]
	Caption=Uppstartsverktyg
	Description=Verktyg som hjälper dig att starta din dator

[devel]
	Caption=Utveckling
	Description=Utvecklingsverktyg så som kompilatorer och assemblerare

[disk]
	Caption=Disk-verktyg
	Description=Verktyg för diskhantering och underhålls

[drivers]
	Caption=Enhetsdrivrutiner
	Description=Drivrutiner för hårdvara och andra enheter

[edit]
	Caption=Redigerare
	Description=Redigerar och enkla ordbehandlare som låter dig redigera textfiler

[emulator]
	Caption=Emulatorer
	Description=Program som emulerar andra system

[games]
	Caption=Spel
	Description=Roliga spel som du kan spela

[gui]
	Caption=Grafiska skrivbord
	Description=Grafiska skrivbordsmiljöer och användargränssnitt

[net]
	Caption=Nätverk
	Description=Verktyg som underlättar nätverkshantering och anslutningar

[sound]
	Caption=Ljudverktyg
	Description=Program för att spela musik- och ljudfiler

[unix]
	Caption=Unix-liknande
	Description=Verktyg som liknar sina motsvarigheter i Unix och Linux

[util]
	Caption=Verktyg
	Description=Generella verktyg och andra användbara progarm som du kan vilja prova

[obsolete]
	Caption=Föråldrade paket
	Description=Pensionerade program som har ersatts med andra program
