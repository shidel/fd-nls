# language: Swedish (Svenska, sv)
# codepage: CP850
# translators: Gemini
# Detta �r en automatiskt genererad text. Om du hittar n�gra fel,
# �r du v�lkommen att korrigera dem och informera FreeDOS-gruppen.

laddad, anv�nder %u bytes.
laddad h�gt, anv�nder %u bytes.
\nKan inte hitta/�ppna Unicode-tabellfil %s!
\nFil %s: Felaktigt inneh�ll eller kan inte l�sas!
inaktiverad.
\n(En annan TSR har tagit Int21 och/eller Int2F)
Inte installerad!
kr�ver minst DOS version 4!
v�xel(ar) godtogs
"
++ FREEWARE ++
Program som st�der l�nga filnamn i ren DOS.
ANV�ND DETTA PROGRAM P� EGEN RISK, DATA F�RLUST �R M�JLIG
�tg�rder:    - (inget)       ladda och/eller aktivera TSR
	     - h eller ?     denna hj�lp
	     - d	     inaktivera DOSLFN
	     - s	     visa status och inst�llningar
?PROFILE
	     - p	     visa profildata
	     - pr	     �terst�ll profildata
	     - pc	     kalibrera profil-timing
?
	     - u	     ladda ur TSR
V�xlar:      - w{+|-}	     * skriv�tkomst
	     - ~{+|-}	     * tilde-anv�ndning (NameNumericTail)
	     - t{+|-}	     * beh�ll l�nga namn (tunneleffekt)
	     - f{+|-}	     * fallback-l�ge: LFN f�r alla enheter
	     - c{+|-}	     * CD-ROM-st�d
	     - i{+|-}	     * �terintr�desl�s (InDOS/RESET)
	     - r{+|-}	     * skrivskydd f�r CD-filer
?USEWINTIME
	     - o[N]	     * st�ll in tidszon N eller l�s TZ
?
	     - z[:|=]tabell  ladda Unicode-tabell (.TBL)
	     - m[:|=]bytes   ange heap-storlek, 600..50000
	     - ms[:|=]bytes  ange kort s�kv�gs-storlek, 16..141
	     - ml[:|=]bytes  ange l�ng s�kv�gs-storlek, 16..1024
	     - mn[:|=]bytes  ange l�ngt namn-storlek, 13..512
	     - p[:|=]s�kv�g  ange arbetskatalog f�r .TBL/.386
Milj�:       LANG=cc	     spr�k f�r meddelanden (NLS\DOSLFN.cc)
?USEWINTIME
	     TZ=xxxNyyy      tidszon N, ingen sommartid
?
Email:	  %s
Download: %s
	  %s
"
aktiv
aktiverad.
borttagen fr�n minnet.
%7lu l�s�tkomster
%7lu skriv�tkomster
%7lu Int21/AH=71-anrop
skriv�tkomst
tilde-anv�ndning
tunneleffekt
CD-ROM-st�d
fallback-l�ge
skrivskyddad bit p� CD-filer
ogiltig heap-storlek
P�
AV
%45s %s\n
katalogen finns inte!
kan inte ange arbetskatalog
kan inte �ndra heap-storlek
v�xel avvisad
 - ladda ur TSR f�rst.
\nDetta program �r oanv�ndbart i en DOS-box i denna Windows-version!
Heap: storlek=%u, anv�nd=%u, ledig=%u, max-tillg�nglig=%u Bytes\n
Anv�ndning av InDOS-flagga och RESET drive
Senaste fel: %u -\s
anv�ndaren nekade skriv�tkomst
kunde inte expandera FAT-katalog
inte tillr�ckligt med minne - �ka heap
kunde inte autoladda Unicode-tabell
?USEWINTIME
Tidszon �r
%45s UTC%+d\n
?
?PROFILE
Profil.\n
Profil �terst�lld.\n
%7lu %2d.%03d %s\n
Kalibrerar profil.\n
Profil-timing-konstant = %lu000\n
Fel vid kalibrering\n
?
