CD.INIT=CD-ROM initiering.
CD.GIVEUP=/p /fLightRed "kan inte l�sa in en l�mplig CD/DVD-drivrutin" /fGrey
CD.ERROR=, /fGrey fel "#%1" - /fLightRed misslyckades /fGrey /p
CD.NO_DRVR= /fGrey kan inte hitta CD-drivrutinen /fYellow "%1" /fGrey - /fLightRed misslyckades /fGrey
CD.TRY_DRVR= /g f�rs�ker att anv�nda CD-drivrutinen /fYellow "%1" /fGrey
CD.TRY_CACHE= /g f�rs�ker att l�sa in /fYellow "%1" /fGrey f�r cachning
CD.TRY_EXT= f�rs�ker att l�sa in CD-till�gget /fYellow "%1" /fGrey
CD.SUCCESS=, /fLightGreen lyckad /fGrey
CD.STATUS=lyckades starta CD-drivrutinen och till�ggen f�r enhet /fLightGreen "%1" /fDarkGrey (%2) /fGrey

CD.DRIVE=CD-ROM konfigurerad som /fLightGreen %1 /fGrey enhet /fDarkGrey (%2) /fGrey
CD.NONE=/fLightRed CD-ROM inte konfigurerad /fGrey

NO_HELP=kan inte hitta hj�lpfil
