# Detta �r den svenska �vers�ttning f�r FreeDOS Password v0.50
#
#               Spr�k: Svenska, sv
#               Kodsida: 850 (Ascii 8bit)
#
# Upphovsman till �vers�ttningen: Sebastian Rasmussen
#
# Alla blanksteg innan text m�ste bevaras och varje rad f�r inte
# inneh�lla n�gra blanksteg p� slutet!
#
0.1:Anv�ndare
0.2:Du m�ste definiera �tminstone en anv�ndare:
0.3:Anv�ndare.:
0.4:L�senord..:
0.5:Anv�ndare
0.6:har lagts till
0.7: VARNING! En fr�mmande person har f�rs�kt att logga in f�rra g�ngen.
0.8:          F�r vidare information, se loggfilen.
0.9: Tryck p� valfri tangent...
0.10:�tkomst nekad!
0.11:Ange anv�ndarnamnet f�r anv�ndaren du vill ta bort:
0.12: Anv�ndare borttagen.
0.13:hittades ej!
0.14:Ange anv�ndaren du vill l�gga till:
0.15:Anv�ndare tillagd
0.16: Anv�ndarnamnet
0.17:anv�nds redan.
0.18: Flaggor:
0.19: /adduser   L�gg till en ny anv�ndare till programmet
0.20: /login     Anv�ndarnamn
0.21: /remuser   Ta bort en anv�ndare fr�n programmet
0.22:har loggat in framg�ngsrikt
0.23:har f�rs�kt att logga in
0.24:har tagits bort
