vpcspkr [hz:][ms]

Generera en ton med hj�lp av den inbyggda h�gtalaren.

    [inga]      Ingen utmatning.
    hz:ms       Anv�nd PC-h�gtalaren f�r att generera en ton med hz frekvens.
                V�nta sedan ms millisekunder. (Ntoera: frekvensen 0 st�nger av
                h�gtalaren. Om ingen frekvens anges antas 0.)
    /D          Detektera metod som anv�nds f�r tidm�tning. (Inte
                kompatibelt med VirtualBox)
    /S          Anv�nd s�ker timer f�r allm�nt bruk. (Standard)
    /I          Anv�nd h�gprecisions timeravbrott. (Inte kompatibelt med
                VirtualBox)

    tba         (Fortfarande under utveckling, mer kommer att annonseras)

