
$OS_NAME$ �r ett DOS-kompatibelt operativsystem med �ppen k�llkod som du kan
anv�nda f�r att spela klassiska DOS-spel, k�ra �ldre aff�rsprogramvara eller
utveckla inbyggda system. Program som fungerar i MS-DOS b�r ocks� k�ra i $OS_NAME$.
*

Du kan spelar dina favorit DOS-spel i $OS_NAME$. Och det finns m�nga bra
klassiska spel att spela: Wolfenstein 3D, Doom, Commander Keen, Rise of the Triad,
Jill of the Jungle, Duke Nukem, och m�nga fler!
*

Beh�ver du �terskapa data fr�n ett gammalt aff�rsprogram? Eller beh�ver du k�ra
en rapport i ditt gamla finanssystem? Bara installera din �ldre programvara under
$OS_NAME$, s� kommer du att klara dig!
*

M�nga inbyggda system k�r p� DOS, �ven om moderna system ist�llet k�r Linux.
Om du underh�ller ett �ldre inbyggt system kanske du k�r DOS. Och $OS_NAME$
passar d� in mycket bra.
*

$OS_NAME$ �r programvara med �ppen k�llkod!
Det kostar ingenting att h�mta och anv�nda $OS_NAME$.
*

FreeDOS Alpha 1 sl�pptes 16:e September 1994. Det �r mer �n 25 �r sedan.
*

Du kan ocks� dela med dig av $OS_NAME$ till andra! Du kan titta p� och redigera
v�r k�llkod eftersom alla $OS_NAME$ program distribueras under licensen GNU
General Public License eller liknande licenser f�r �ppen k�lkod.
*

$OS_NAME$ har alltid handlat om att utvecklare samlas f�r att skriva kod.
Bes�k $OS_NAME$-projektets webbplats f�r vidare information om hur du kan
bidra till $OS_NAME$.
*

Har du fr�gor om hur du st�ller in eller anv�nder $OS_NAME$? Kolla p�
s�ndlistan f�r FreeDOS-anv�ndare p� webbplatsens Forumsida.
