AUTO_DONE=Behandling av uppstartsfiler klar /fCyan %1 /a7 och /fCyan %2 /a7
AUTO_HELP=Skriv /fWhite %1 /fGray f�r att f� hj�lp med kommandon och navigering.
AUTO_WELCOME=V�lkommen till operativsystemet /fGreen %1 /fCyan %2 /fGray ( /s- /fYellow "%3" /fGray )
