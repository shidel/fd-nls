version
Detta verktyg kan utv�rdera ett givet matematiskt uttryck
Skrivet av Laaca under GNU/GPL-licensen.
Anv�nd vanlig notation f�r datorer. Upph�jningar anges med "^"-operatorn.
Ange ett matematiskt uttryck:
Dessa funktioner st�ds
Du kan ocks� anv�nda dessa bitoperatorer: AND, OR, XOR
fel vid pos. n.
division med noll
ogiltigt argument i rot
flyttalsargument i bitoperation
f�r stort resultat i matteoperation
f�r litet resultat i matteoperation
noll eller negativ logaritm


# swedish, sv, cp850/858
