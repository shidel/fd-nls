vpause [flaggor]

Enkel v�ntan p� tangenttryckning eller tidsgr�ns.

    [inga]      V�nta f�r evigt p� en tangenttryckning.
    (/T)        F�r�ldrad. Numera, /D.
    /D sekunder F�rdr�jing i sekunder att v�nta innan pausens tidgr�ns l�per
                ut. (returnerar errorlevel 1)
    CTRL-C      N�r angivet och Ctrl-C trycks, avsluta med errorlevel 200.

    tba         (Fortfarande under utveckling, mer kommer att annonseras)

