[repository]

	Caption=FreeDOS 1.3 nedladdningar
	Description=Programvaruförråd för hämtningar och uppdateringar för FreeDOS 1.3
